library verilog;
use verilog.vl_types.all;
entity TestClockDivider is
end TestClockDivider;
