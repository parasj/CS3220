module Controller(in, src_index1, src_index2, dst_index, alu_op, imm, cmd_flag);

endmodule