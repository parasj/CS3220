module ClockDivider (
	inclk0,
	c0,
	locked);

	input	  inclk0;
	output	  c0;
	output	  locked; // clock is paused when locked is 1

  // Implement this yourself
  // Slow down the clock to ensure the cycle is long enough for all operations to execute
  // If you don't, you might get weird errors
  

endmodule
