module Controller(in, src_index1, src_index2, dst_index, imm, alu_op, alu_mux, dstdata_mux, reg_wrt_en, mem_wrt_en, nextpc_mux, cmd_flag);
	input [31:0] in;
	input cmd_flag;
	output[3:0] src_index1, src_index2, dst_index;
	output[1:0] alu_mux, dstdata_mux, nextpc_mux;
	output reg_wrt_en, mem_wrt_en;
	output[4:0] alu_op;
	output[15:0] imm;

	wire [3:0] op;
	wire [3:0] fn;
	wire [8:0] x;
	wire [12:0] out;

	assign src_index1 = in[19:16];
	assign src_index2 = in[15:12];
	assign dst_index = in[23:20];
	assign imm = in[15:0];
	assign x = {in[31:24], cmd_flag};
	assign alu_op = out[12:8];
	assign alu_mux = out[7:6];
	assign dstdata_mux = out[5:4];
	assign reg_wrt_en = out[3];
	assign mem_wrt_en = out[2];
	assign nextpc_mux = out[1:0];

	assign out =	(x == 9'b110001110) ? 13'b0000100001000 :
					(x == 9'b110001100) ? 13'b0001000001000 :
					(x == 9'b110000000) ? 13'b0001100001000 :
					(x == 9'b110000010) ? 13'b0010000001000 :
					(x == 9'b110000100) ? 13'b0010100001000 :
					(x == 9'b110010000) ? 13'b0011000001000 :
					(x == 9'b110010010) ? 13'b0011100001000 :
					(x == 9'b110010100) ? 13'b0100000001000 :
					(x == 9'b010001110) ? 13'b0000101001000 :
					(x == 9'b010001100) ? 13'b0001001001000 :
					(x == 9'b010000000) ? 13'b0001101001000 :
					(x == 9'b010000010) ? 13'b0010001001000 :
					(x == 9'b010000100) ? 13'b0010101001000 :
					(x == 9'b010010000) ? 13'b0011001001000 :
					(x == 9'b010010010) ? 13'b0011101001000 :
					(x == 9'b010010100) ? 13'b0100001001000 :
					(x == 9'b010011110) ? 13'b0100101001000 :
					(x == 9'b011100000) ? 13'b0000100101000 :
					(x == 9'b001100000) ? 13'b0000100010100 :
					(x == 9'b110100110) ? 13'b0101000001000 :
					(x == 9'b110101100) ? 13'b0101100001000 :
					(x == 9'b110110010) ? 13'b0110000001000 :
					(x == 9'b110111000) ? 13'b0110100001000 :
					(x == 9'b110100000) ? 13'b0111000001000 :
					(x == 9'b110101010) ? 13'b0111100001000 :
					(x == 9'b110110100) ? 13'b1000000001000 :
					(x == 9'b110111110) ? 13'b1000100001000 :
					(x == 9'b010100110) ? 13'b0101001001000 :
					(x == 9'b010101100) ? 13'b0101101001000 :
					(x == 9'b010110010) ? 13'b0110001001000 :
					(x == 9'b010111000) ? 13'b0110101001000 :
					(x == 9'b010100000) ? 13'b0111001001000 :
					(x == 9'b010101010) ? 13'b0111101001000 :
					(x == 9'b010110100) ? 13'b1000001001000 :
					(x == 9'b010111110) ? 13'b1000101001000 :
					(x == 9'b001000110) ? 13'b0101000000000 :
					(x == 9'b001001100) ? 13'b0101100000000 :
					(x == 9'b001010010) ? 13'b0110000000000 :
					(x == 9'b001011000) ? 13'b0110100000000 :
					(x == 9'b001000100) ? 13'b1001000000000 :
					(x == 9'b001011010) ? 13'b1001100000000 :
					(x == 9'b001010000) ? 13'b1010000000000 :
					(x == 9'b001000000) ? 13'b0111000000000 :
					(x == 9'b001001010) ? 13'b0111100000000 :
					(x == 9'b001010100) ? 13'b1000000000000 :
					(x == 9'b001010110) ? 13'b1000100000000 :
					(x == 9'b001000010) ? 13'b1010100000000 :
					(x == 9'b001011100) ? 13'b1011000000000 :
					(x == 9'b001011110) ? 13'b1011100000000 :
					(x == 9'b011000000) ? 13'b0000110101000 :
					(x == 9'b110001111) ? 13'b0000100001000 :
					(x == 9'b110001101) ? 13'b0001000001000 :
					(x == 9'b110000001) ? 13'b0001100001000 :
					(x == 9'b110000011) ? 13'b0010000001000 :
					(x == 9'b110000101) ? 13'b0010100001000 :
					(x == 9'b110010001) ? 13'b0011000001000 :
					(x == 9'b110010011) ? 13'b0011100001000 :
					(x == 9'b110010101) ? 13'b0100000001000 :
					(x == 9'b010001111) ? 13'b0000101001000 :
					(x == 9'b010001101) ? 13'b0001001001000 :
					(x == 9'b010000001) ? 13'b0001101001000 :
					(x == 9'b010000011) ? 13'b0010001001000 :
					(x == 9'b010000101) ? 13'b0010101001000 :
					(x == 9'b010010001) ? 13'b0011001001000 :
					(x == 9'b010010011) ? 13'b0011101001000 :
					(x == 9'b010010101) ? 13'b0100001001000 :
					(x == 9'b010011111) ? 13'b0100101001000 :
					(x == 9'b011100001) ? 13'b0000100101000 :
					(x == 9'b001100001) ? 13'b0000100010100 :
					(x == 9'b110100111) ? 13'b0101000001000 :
					(x == 9'b110101101) ? 13'b0101100001000 :
					(x == 9'b110110011) ? 13'b0110000001000 :
					(x == 9'b110111001) ? 13'b0110100001000 :
					(x == 9'b110100001) ? 13'b0111000001000 :
					(x == 9'b110101011) ? 13'b0111100001000 :
					(x == 9'b110110101) ? 13'b1000000001000 :
					(x == 9'b110111111) ? 13'b1000100001000 :
					(x == 9'b010100111) ? 13'b0101001001000 :
					(x == 9'b010101101) ? 13'b0101101001000 :
					(x == 9'b010110011) ? 13'b0110001001000 :
					(x == 9'b010111001) ? 13'b0110101001000 :
					(x == 9'b010100001) ? 13'b0111001001000 :
					(x == 9'b010101011) ? 13'b0111101001000 :
					(x == 9'b010110101) ? 13'b1000001001000 :
					(x == 9'b010111111) ? 13'b1000101001000 :
					(x == 9'b001000111) ? 13'b0101000000001 :
					(x == 9'b001001101) ? 13'b0101100000001 :
					(x == 9'b001010011) ? 13'b0110000000001 :
					(x == 9'b001011001) ? 13'b0110100000001 :
					(x == 9'b001000101) ? 13'b1001000000001 :
					(x == 9'b001011011) ? 13'b1001100000001 :
					(x == 9'b001010001) ? 13'b1010000000001 :
					(x == 9'b001000001) ? 13'b0111000000001 :
					(x == 9'b001001011) ? 13'b0111100000001 :
					(x == 9'b001010101) ? 13'b1000000000001 :
					(x == 9'b001010111) ? 13'b1000100000001 :
					(x == 9'b001000011) ? 13'b1010100000001 :
					(x == 9'b001011101) ? 13'b1011000000001 :
					(x == 9'b001011111) ? 13'b1011100000001 :
					(x == 9'b011000001) ? 13'b0000110101010 :
					{13{x}};
endmodule