library verilog;
use verilog.vl_types.all;
entity Timer is
    port(
        SW              : in     vl_logic_vector(7 downto 0);
        KEY             : in     vl_logic_vector(2 downto 0);
        LEDR            : out    vl_logic_vector(9 downto 0);
        HEX0            : out    vl_logic_vector(6 downto 0);
        HEX1            : out    vl_logic_vector(6 downto 0);
        HEX2            : out    vl_logic_vector(6 downto 0);
        HEX3            : out    vl_logic_vector(6 downto 0);
        CLOCK_50        : in     vl_logic
    );
end Timer;
