module MEM_WB_Buffer(clk, reset, en, reg_file_wrt_en_in, reg_file_wrt_en_out, dst_ind_in,
	dst_ind_out, end_res_in, end_res_out);

endmodule