module DummyMemory2(addr, dataOut);
	parameter MEM_INIT_FILE;
	parameter ADDR_BIT_WIDTH = 11;
	parameter DATA_BIT_WIDTH = 32;
	parameter N_WORDS = (1 << ADDR_BIT_WIDTH);
	
	input[ADDR_BIT_WIDTH - 1: 0] addr;
	output[DATA_BIT_WIDTH - 1: 0] dataOut;

	reg[DATA_BIT_WIDTH - 1: 0] data[0: N_WORDS - 1];
	
	assign dataOut = data[addr];

	initial begin
		data[16] = 32'h4fe00000;
		data[17] = 32'h47ee2000;
		data[18] = 32'h4fc0f000;
		data[19] = 32'h40660000;
		data[20] = 32'h306c0004;
		data[21] = 32'h47460100;
		data[22] = 32'h47541000;
		data[23] = 32'h47760009;
		data[24] = 32'h30740000;
		data[25] = 32'h4777000d;
		data[26] = 32'h47440004;
		data[27] = 32'h2545fffc;
		data[28] = 32'h60f6002d;
		data[29] = 32'h4776012c;
		data[30] = 32'h307c0000;
		data[31] = 32'h47060100;
		data[32] = 32'h47101000;
		data[33] = 32'h60f60055;
		data[34] = 32'h60f6003a;
		data[35] = 32'h47060100;
		data[36] = 32'h47101000;
		data[37] = 32'h60f60047;
		data[38] = 32'h60f6002d;
		data[39] = 32'h4777ffff;
		data[40] = 32'h307c0000;
		data[41] = 32'h2170fff5;
		data[42] = 32'hc8466000;
		data[43] = 32'h306c0004;
		data[44] = 32'h2046fffd;
		data[45] = 32'h47060100;
		data[46] = 32'h47101000;
		data[47] = 32'h47260009;
		data[48] = 32'h70400000;
		data[49] = 32'h26420004;
		data[50] = 32'h304c0000;
		data[51] = 32'h475603e0;
		data[52] = 32'h305c0004;
		data[53] = 32'h2044fffc;
		data[54] = 32'h4722000d;
		data[55] = 32'h47000004;
		data[56] = 32'h2501fff7;
		data[57] = 32'h609f0000;
		data[58] = 32'h47160100;
		data[59] = 32'h47011000;
		data[60] = 32'h47260009;
		data[61] = 32'h46000004;
		data[62] = 32'h70500000;
		data[63] = 32'h26250004;
		data[64] = 32'h305c0000;
		data[65] = 32'h4746001f;
		data[66] = 32'h304c0004;
		data[67] = 32'h2054fffc;
		data[68] = 32'h4722000d;
		data[69] = 32'h2510fff7;
		data[70] = 32'h609f0000;
		data[71] = 32'h2601000c;
		data[72] = 32'h70400000;
		data[73] = 32'h47200004;
		data[74] = 32'h26210006;
		data[75] = 32'h70520000;
		data[76] = 32'h2c450002;
		data[77] = 32'h30420000;
		data[78] = 32'hc7456000;
		data[79] = 32'h47220004;
		data[80] = 32'h2045fff9;
		data[81] = 32'h30400000;
		data[82] = 32'h47000004;
		data[83] = 32'h2001fff3;
		data[84] = 32'h609f0000;
		data[85] = 32'h47400000;
		data[86] = 32'h2641000b;
		data[87] = 32'h47540004;
		data[88] = 32'h26510007;
		data[89] = 32'h70240000;
		data[90] = 32'h70350000;
		data[91] = 32'h2a230002;
		data[92] = 32'h30250000;
		data[93] = 32'h30340000;
		data[94] = 32'h47550004;
		data[95] = 32'h2000fff8;
		data[96] = 32'h47440004;
	end
endmodule