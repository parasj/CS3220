library verilog;
use verilog.vl_types.all;
entity TestAdderSubtractor is
end TestAdderSubtractor;
