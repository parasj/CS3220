library verilog;
use verilog.vl_types.all;
entity TestClockMultipler is
end TestClockMultipler;
