module DEC_EXE_Buffer(clk, reset, en, pc_in, pc_out, src1_in, src1_out, src2_in, src2_out, imm_in, imm_out, alu_mux_op);
	parameter BIT_WIDTH = 32;
	parameter INST_BIT_WIDTH				 = 32;
	parameter REG_INDEX_BIT_WIDTH 		 = 4;

	input clk, reset, en;
	
endmodule