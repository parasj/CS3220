module Controller(in, src_index1, src_index2, dst_index, imm, alu_op, alu_mux, dstdata_mux, reg_wrt_en, mem_wrt_en, nextpc_mux, cmd_flag, fn_exe_in, fn_exe_out);
	parameter INST_BIT_WIDTH = 32;
	input [INST_BIT_WIDTH - 1 : 0] in;
	
	input cmd_flag;
	output[3:0] src_index1, src_index2, dst_index;
	output alu_mux, dstdata_mux, nextpc_mux;
	output reg_wrt_en, mem_wrt_en;
	output [4:0] alu_op;
	output[15:0] imm;
	input[3:0] fn_exe_in;
	input[3:0] fn_exe_out;

	wire [3:0] op;
	wire [3:0] fn;
	wire [8:0] x;
	wire [8:0] out;
	assign fn = in[31:28];
	assign src_index1 = (fn == 4'b0010) ? in[23:20] : in[19:16];
	assign src_index2 = (fn == 4'b0010) ? in[19:16] : (fn == 4'b0011) ? in [23:20] : in[15:12];
	assign dst_index = in[23:20];
	assign imm = (fn == 4'b0110) ? in[15:0] << 2 : in[15:0];
	assign x = {in[INST_BIT_WIDTH - 1 : 24]};
	assign alu_op = out[8:4];
	assign alu_mux = out[3];
	assign dstdata_mux = out[2];
	assign reg_wrt_en = out[1];
	assign mem_wrt_en = out[0];
	assign fn_exe_out = fn;

	assign nextpc_mux =	(cmd_flag == 1 & (fn_exe_in == 4'b0110 | fn_exe_in == 4'b0010)) ? 1 : 0;

	assign out =	(x == 8'b11000111) ? 9'b000010010 :
					(x == 8'b11000110) ? 9'b000100010 :
					(x == 8'b11000000) ? 9'b000110010 :
					(x == 8'b11000001) ? 9'b001000010 :
					(x == 8'b11000010) ? 9'b001010010 :
					(x == 8'b11001000) ? 9'b001100010 :
					(x == 8'b11001001) ? 9'b001110010 :
					(x == 8'b11001010) ? 9'b010000010 :
					(x == 8'b01000111) ? 9'b000011010 :
					(x == 8'b01000110) ? 9'b000101010 :
					(x == 8'b01000000) ? 9'b000111010 :
					(x == 8'b01000001) ? 9'b001001010 :
					(x == 8'b01000010) ? 9'b001011010 :
					(x == 8'b01001000) ? 9'b001101010 :
					(x == 8'b01001001) ? 9'b001111010 :
					(x == 8'b01001010) ? 9'b010001010 :
					(x == 8'b01001111) ? 9'b010011010 :
					(x == 8'b01110000) ? 9'b000011110 :
					(x == 8'b00110000) ? 9'b000011001 :
					(x == 8'b11010011) ? 9'b010100010 :
					(x == 8'b11010110) ? 9'b010110010 :
					(x == 8'b11011001) ? 9'b011000010 :
					(x == 8'b11011100) ? 9'b011010010 :
					(x == 8'b11010000) ? 9'b011100010 :
					(x == 8'b11010101) ? 9'b011110010 :
					(x == 8'b11011010) ? 9'b100000010 :
					(x == 8'b11011111) ? 9'b100010010 :
					(x == 8'b01010011) ? 9'b010101010 :
					(x == 8'b01010110) ? 9'b010111010 :
					(x == 8'b01011001) ? 9'b011001010 :
					(x == 8'b01011100) ? 9'b011011010 :
					(x == 8'b01010000) ? 9'b011101010 :
					(x == 8'b01010101) ? 9'b011111010 :
					(x == 8'b01011010) ? 9'b100001010 :
					(x == 8'b01011111) ? 9'b100011010 :
					(x == 8'b00100011) ? 9'b010100000 :
					(x == 8'b00100110) ? 9'b010110000 :
					(x == 8'b00101001) ? 9'b011000000 :
					(x == 8'b00101100) ? 9'b011010000 :
					(x == 8'b00100010) ? 9'b100100000 :
					(x == 8'b00101101) ? 9'b100110000 :
					(x == 8'b00101000) ? 9'b101000000 :
					(x == 8'b00100000) ? 9'b011100000 :
					(x == 8'b00100101) ? 9'b011110000 :
					(x == 8'b00101010) ? 9'b100000000 :
					(x == 8'b00101011) ? 9'b100010000 :
					(x == 8'b00100001) ? 9'b101010000 :
					(x == 8'b00101110) ? 9'b101100000 :
					(x == 8'b00101111) ? 9'b101110000 :
					(x == 8'b01100000) ? 9'b000011110 :
					(x == 8'b11000111) ? 9'b000010010 :
					(x == 8'b11000110) ? 9'b000100010 :
					(x == 8'b11000000) ? 9'b000110010 :
					(x == 8'b11000001) ? 9'b001000010 :
					(x == 8'b11000010) ? 9'b001010010 :
					(x == 8'b11001000) ? 9'b001100010 :
					(x == 8'b11001001) ? 9'b001110010 :
					(x == 8'b11001010) ? 9'b010000010 :
					(x == 8'b01000111) ? 9'b000011010 :
					(x == 8'b01000110) ? 9'b000101010 :
					(x == 8'b01000000) ? 9'b000111010 :
					(x == 8'b01000001) ? 9'b001001010 :
					(x == 8'b01000010) ? 9'b001011010 :
					(x == 8'b01001000) ? 9'b001101010 :
					(x == 8'b01001001) ? 9'b001111010 :
					(x == 8'b01001010) ? 9'b010001010 :
					(x == 8'b01001111) ? 9'b010011010 :
					(x == 8'b01110000) ? 9'b000011110 :
					(x == 8'b00110000) ? 9'b000011001 :
					(x == 8'b11010011) ? 9'b010100010 :
					(x == 8'b11010110) ? 9'b010110010 :
					(x == 8'b11011001) ? 9'b011000010 :
					(x == 8'b11011100) ? 9'b011010010 :
					(x == 8'b11010000) ? 9'b011100010 :
					(x == 8'b11010101) ? 9'b011110010 :
					(x == 8'b11011010) ? 9'b100000010 :
					(x == 8'b11011111) ? 9'b100010010 :
					(x == 8'b01010011) ? 9'b010101010 :
					(x == 8'b01010110) ? 9'b010111010 :
					(x == 8'b01011001) ? 9'b011001010 :
					(x == 8'b01011100) ? 9'b011011010 :
					(x == 8'b01010000) ? 9'b011101010 :
					(x == 8'b01010101) ? 9'b011111010 :
					(x == 8'b01011010) ? 9'b100001010 :
					(x == 8'b01011111) ? 9'b100011010 :
					(x == 8'b00100011) ? 9'b010100000 :
					(x == 8'b00100110) ? 9'b010110000 :
					(x == 8'b00101001) ? 9'b011000000 :
					(x == 8'b00101100) ? 9'b011010000 :
					(x == 8'b00100010) ? 9'b100100000 :
					(x == 8'b00101101) ? 9'b100110000 :
					(x == 8'b00101000) ? 9'b101000000 :
					(x == 8'b00100000) ? 9'b011100000 :
					(x == 8'b00100101) ? 9'b011110000 :
					(x == 8'b00101010) ? 9'b100000000 :
					(x == 8'b00101011) ? 9'b100010000 :
					(x == 8'b00100001) ? 9'b101010000 :
					(x == 8'b00101110) ? 9'b101100000 :
					(x == 8'b00101111) ? 9'b101110000 :
					(x == 8'b01100000) ? 9'b000011110 :
					{13{x}};
endmodule