module TestClockMultipler;
	
endmodule