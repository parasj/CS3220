module TestClockMultipler;
	ClockMultiplier()
end