module DummyMemory(addr, dataOut);
	parameter MEM_INIT_FILE;
	parameter ADDR_BIT_WIDTH = 11;
	parameter DATA_BIT_WIDTH = 32;
	parameter N_WORDS = (1 << ADDR_BIT_WIDTH);
	
	input[ADDR_BIT_WIDTH - 1: 0] addr;
	output[DATA_BIT_WIDTH - 1: 0] dataOut;

	reg[DATA_BIT_WIDTH - 1: 0] data[0: N_WORDS - 1];
	
	assign dataOut = data[addr];

	initial begin
		data[0] = 32'h20440008;
		data[1] = 32'h47770001;
		data[2] = 32'h47770001;
		data[3] = 32'h47770001;
		data[4] = 32'h47770001;
		data[5] = 32'h47770001;
		data[6] = 32'h47770001;
		data[7] = 32'h47770001;
		data[8] = 32'h47770001;
		data[9] = 32'h4fc0f000;
		data[10] = 32'h40660000;
		data[11] = 32'hc8466000;
		data[12] = 32'h304c0004;
		data[13] = 32'h47460bad;
		data[14] = 32'h304c0000;
		data[16] = 32'h47860bef;
		data[17] = 32'hc2ddd000;
		data[18] = 32'h4fc0f000;
		data[19] = 32'h4f600000;
		data[20] = 32'h47660001;
		data[21] = 32'h306c0004;
		data[22] = 32'h47660001;
		data[23] = 32'h306c0004;
		data[24] = 32'h474dffff;
		data[25] = 32'h475d0002;
		data[26] = 32'h470d0001;
		data[27] = 32'hc7145000;
		data[28] = 32'h26010004;
		data[29] = 32'hc84dd000;
		data[30] = 32'h304c0004;
		data[31] = 32'h300c0000;
		data[32] = 32'h2044fffc;
		data[33] = 32'h47660001;
		data[34] = 32'h306c0004;
		data[35] = 32'h474d0007;
		data[36] = 32'h47540003;
		data[37] = 32'hc7055000;
		data[38] = 32'h41100025;
		data[39] = 32'h402100d1;
		data[40] = 32'hc2001000;
		data[41] = 32'hc1104000;
		data[42] = 32'hc9242000;
		data[43] = 32'hc8321000;
		data[44] = 32'hc6142000;
		data[45] = 32'hc0412000;
		data[46] = 32'hca114000;
		data[47] = 32'hc2223000;
		data[48] = 32'hc6002000;
		data[49] = 32'hc7010000;
		data[50] = 32'h475dfff8;
		data[51] = 32'h25050004;
		data[52] = 32'hc84dd000;
		data[53] = 32'h304c0004;
		data[54] = 32'h300c0000;
		data[55] = 32'h2044fffc;
		data[56] = 32'h47660001;
		data[57] = 32'h306c0004;
		data[58] = 32'h471d0001;
		data[59] = 32'h474d004b;
		data[60] = 32'h475d0022;
		data[61] = 32'h470dffb0;
		data[62] = 32'hdc245000;
		data[63] = 32'h252d0045;
		data[64] = 32'h47660001;
		data[65] = 32'h306c0004;
		data[66] = 32'hd9245000;
		data[67] = 32'h252d0041;
		data[68] = 32'h47660001;
		data[69] = 32'h306c0004;
		data[70] = 32'hd6245000;
		data[71] = 32'h252d003d;
		data[72] = 32'h47660001;
		data[73] = 32'h306c0004;
		data[74] = 32'hd5245000;
		data[75] = 32'h25210039;
		data[76] = 32'h47660001;
		data[77] = 32'h306c0004;
		data[78] = 32'hdf245000;
		data[79] = 32'h25210035;
		data[80] = 32'h47660001;
		data[81] = 32'h306c0004;
		data[82] = 32'hda245000;
		data[83] = 32'h25210031;
		data[84] = 32'h47660001;
		data[85] = 32'h306c0004;
		data[86] = 32'hdc255000;
		data[87] = 32'h2521002d;
		data[88] = 32'h47660001;
		data[89] = 32'h306c0004;
		data[90] = 32'hd9255000;
		data[91] = 32'h252d0029;
		data[92] = 32'h47660001;
		data[93] = 32'h306c0004;
		data[94] = 32'hd6255000;
		data[95] = 32'h25210025;
		data[96] = 32'h47660001;
		data[97] = 32'h306c0004;
		data[98] = 32'hd5255000;
		data[99] = 32'h252d0021;
		data[100] = 32'h47660001;
		data[101] = 32'h306c0004;
		data[102] = 32'hdf255000;
		data[103] = 32'h252d001d;
		data[104] = 32'h47660001;
		data[105] = 32'h306c0004;
		data[106] = 32'hda255000;
		data[107] = 32'h25210019;
		data[108] = 32'h47660001;
		data[109] = 32'h306c0004;
		data[110] = 32'hdc204000;
		data[111] = 32'h25210015;
		data[112] = 32'h47660001;
		data[113] = 32'h306c0004;
		data[114] = 32'hd9204000;
		data[115] = 32'h25210011;
		data[116] = 32'h47660001;
		data[117] = 32'h306c0004;
		data[118] = 32'hd6204000;
		data[119] = 32'h252d000d;
		data[120] = 32'h47660001;
		data[121] = 32'h306c0004;
		data[122] = 32'hd5204000;
		data[123] = 32'h25210009;
		data[124] = 32'h47660001;
		data[125] = 32'h306c0004;
		data[126] = 32'hdf204000;
		data[127] = 32'h252d0005;
		data[128] = 32'h47660001;
		data[129] = 32'h306c0004;
		data[130] = 32'hda204000;
		data[131] = 32'h252d0001;
		data[132] = 32'h20440004;
		data[133] = 32'hc84cc000;
		data[134] = 32'h304c0004;
		data[135] = 32'h302c0000;
		data[136] = 32'h2044fffc;
		data[137] = 32'h47660001;
		data[138] = 32'h306c0004;
		data[139] = 32'h474d0037;
		data[140] = 32'h475d00e1;
		data[141] = 32'h472d0400;
		data[142] = 32'h30420000;
		data[143] = 32'h30520004;
		data[144] = 32'h47220004;
		data[145] = 32'h70020000;
		data[146] = 32'h25050002;
		data[147] = 32'h7002fffc;
		data[148] = 32'h26040004;
		data[149] = 32'hc84dd000;
		data[150] = 32'h304c0004;
		data[151] = 32'h300c0000;
		data[152] = 32'h2044fffc;
		data[153] = 32'h47660001;
		data[154] = 32'h306c0004;
		data[155] = 32'h475d009f;
		data[156] = 32'hc7555000;
		data[157] = 32'hc7555000;
		data[158] = 32'h604d00a0;
		data[159] = 32'h20440006;
		data[160] = 32'h25450001;
		data[161] = 32'h60540000;
		data[162] = 32'hc84dd000;
		data[163] = 32'h304c0004;
		data[164] = 32'h304c0000;
		data[165] = 32'h2044fffc;
		data[166] = 32'h47660001;
		data[167] = 32'h306c0004;
		data[168] = 32'h705c0010;
		data[169] = 32'h305c0000;
		data[170] = 32'h265dfffd;
		data[171] = 32'h705c0010;
		data[172] = 32'h305c0000;
		data[173] = 32'h255dfffd;
		data[174] = 32'hc84dd000;
		data[175] = 32'h304c0004;
		data[176] = 32'h304c0000;
		data[177] = 32'h2044fffc;
	end
endmodule