module Processor(SW, KEY, LEDR, HEX0, HEX1, HEX2, HEX3, CLOCK_50);
	input	[9:0] SW;
	input	[3:0] KEY;
	input	CLOCK_50;
	output	[9:0] LEDR;
	output	[6:0] HEX0, HEX1, HEX2, HEX3;

	
endmodule